-- Effect_Pedal_Memory_Controller.vhd

-- Generated using ACDS version 20.1 720

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Effect_Pedal_Memory_Controller is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity Effect_Pedal_Memory_Controller;

architecture rtl of Effect_Pedal_Memory_Controller is
	component Effect_Pedal_Memory_Controller_SDRAMtest_0 is
		port (
			Avalon_Pipelined_MM_0_avm_m0_address       : in    std_logic_vector(25 downto 0) := (others => 'X'); -- address
			Avalon_Pipelined_MM_0_avm_m0_read          : in    std_logic                     := 'X';             -- read
			Avalon_Pipelined_MM_0_avm_m0_waitrequest   : out   std_logic;                                        -- waitrequest
			Avalon_Pipelined_MM_0_avm_m0_readdata      : out   std_logic_vector(31 downto 0);                    -- readdata
			Avalon_Pipelined_MM_0_avm_m0_readdatavalid : out   std_logic;                                        -- readdatavalid
			Avalon_Pipelined_MM_0_avm_m0_write         : in    std_logic                     := 'X';             -- write
			Avalon_Pipelined_MM_0_avm_m0_writedata     : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			Avalon_Pipelined_MM_0_reset_reset          : out   std_logic;                                        -- reset
			de10_clk_clk                               : in    std_logic                     := 'X';             -- clk
			reset_reset_n                              : in    std_logic                     := 'X';             -- reset_n
			sdram_clk_clk                              : out   std_logic;                                        -- clk
			sdram_wire_addr                            : out   std_logic_vector(12 downto 0);                    -- addr
			sdram_wire_ba                              : out   std_logic_vector(1 downto 0);                     -- ba
			sdram_wire_cas_n                           : out   std_logic;                                        -- cas_n
			sdram_wire_cke                             : out   std_logic;                                        -- cke
			sdram_wire_cs_n                            : out   std_logic;                                        -- cs_n
			sdram_wire_dq                              : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			sdram_wire_dqm                             : out   std_logic_vector(1 downto 0);                     -- dqm
			sdram_wire_ras_n                           : out   std_logic;                                        -- ras_n
			sdram_wire_we_n                            : out   std_logic                                         -- we_n
		);
	end component Effect_Pedal_Memory_Controller_SDRAMtest_0;

begin

	sdramtest_0 : component Effect_Pedal_Memory_Controller_SDRAMtest_0
		port map (
			Avalon_Pipelined_MM_0_avm_m0_address       => open,          -- Avalon_Pipelined_MM_0_avm_m0.address
			Avalon_Pipelined_MM_0_avm_m0_read          => open,          --                             .read
			Avalon_Pipelined_MM_0_avm_m0_waitrequest   => open,          --                             .waitrequest
			Avalon_Pipelined_MM_0_avm_m0_readdata      => open,          --                             .readdata
			Avalon_Pipelined_MM_0_avm_m0_readdatavalid => open,          --                             .readdatavalid
			Avalon_Pipelined_MM_0_avm_m0_write         => open,          --                             .write
			Avalon_Pipelined_MM_0_avm_m0_writedata     => open,          --                             .writedata
			Avalon_Pipelined_MM_0_reset_reset          => open,          --  Avalon_Pipelined_MM_0_reset.reset
			de10_clk_clk                               => clk_clk,       --                     de10_clk.clk
			reset_reset_n                              => reset_reset_n, --                        reset.reset_n
			sdram_clk_clk                              => open,          --                    sdram_clk.clk
			sdram_wire_addr                            => open,          --                   sdram_wire.addr
			sdram_wire_ba                              => open,          --                             .ba
			sdram_wire_cas_n                           => open,          --                             .cas_n
			sdram_wire_cke                             => open,          --                             .cke
			sdram_wire_cs_n                            => open,          --                             .cs_n
			sdram_wire_dq                              => open,          --                             .dq
			sdram_wire_dqm                             => open,          --                             .dqm
			sdram_wire_ras_n                           => open,          --                             .ras_n
			sdram_wire_we_n                            => open           --                             .we_n
		);

end architecture rtl; -- of Effect_Pedal_Memory_Controller
