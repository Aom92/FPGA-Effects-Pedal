// ADC.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module ADC (
		input  wire        adc_command_valid,          //  adc_command.valid
		input  wire [4:0]  adc_command_channel,        //             .channel
		input  wire        adc_command_startofpacket,  //             .startofpacket
		input  wire        adc_command_endofpacket,    //             .endofpacket
		output wire        adc_command_ready,          //             .ready
		output wire        adc_response_valid,         // adc_response.valid
		output wire        adc_response_startofpacket, //             .startofpacket
		output wire        adc_response_endofpacket,   //             .endofpacket
		output wire [0:0]  adc_response_empty,         //             .empty
		output wire [4:0]  adc_response_channel,       //             .channel
		output wire [11:0] adc_response_data,          //             .data
		input  wire        clk_adc_clk,                //      clk_adc.clk
		input  wire        reset_reset_n               //        reset.reset_n
	);

	wire    altpll_0_c0_clk;                // altpll_0:c0 -> modular_adc_0:adc_pll_clock_clk
	wire    altpll_0_locked_conduit_export; // altpll_0:locked -> modular_adc_0:adc_pll_locked_export
	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> [altpll_0:reset, modular_adc_0:reset_sink_reset_n]

	ADC_altpll_0 altpll_0 (
		.clk                (clk_adc_clk),                    //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset), // inclk_interface_reset.reset
		.read               (),                               //             pll_slave.read
		.write              (),                               //                      .write
		.address            (),                               //                      .address
		.readdata           (),                               //                      .readdata
		.writedata          (),                               //                      .writedata
		.c0                 (altpll_0_c0_clk),                //                    c0.clk
		.locked             (altpll_0_locked_conduit_export), //        locked_conduit.export
		.scandone           (),                               //           (terminated)
		.scandataout        (),                               //           (terminated)
		.c1                 (),                               //           (terminated)
		.c2                 (),                               //           (terminated)
		.c3                 (),                               //           (terminated)
		.c4                 (),                               //           (terminated)
		.areset             (1'b0),                           //           (terminated)
		.phasedone          (),                               //           (terminated)
		.phasecounterselect (3'b000),                         //           (terminated)
		.phaseupdown        (1'b0),                           //           (terminated)
		.phasestep          (1'b0),                           //           (terminated)
		.scanclk            (1'b0),                           //           (terminated)
		.scanclkena         (1'b0),                           //           (terminated)
		.scandata           (1'b0),                           //           (terminated)
		.configupdate       (1'b0)                            //           (terminated)
	);

	ADC_modular_adc_0 #(
		.is_this_first_or_second_adc (1)
	) modular_adc_0 (
		.clock_clk              (clk_adc_clk),                     //          clock.clk
		.reset_sink_reset_n     (~rst_controller_reset_out_reset), //     reset_sink.reset_n
		.adc_pll_clock_clk      (altpll_0_c0_clk),                 //  adc_pll_clock.clk
		.adc_pll_locked_export  (altpll_0_locked_conduit_export),  // adc_pll_locked.export
		.command_valid          (adc_command_valid),               //        command.valid
		.command_channel        (adc_command_channel),             //               .channel
		.command_startofpacket  (adc_command_startofpacket),       //               .startofpacket
		.command_endofpacket    (adc_command_endofpacket),         //               .endofpacket
		.command_ready          (adc_command_ready),               //               .ready
		.response_valid         (adc_response_valid),              //       response.valid
		.response_startofpacket (adc_response_startofpacket),      //               .startofpacket
		.response_endofpacket   (adc_response_endofpacket),        //               .endofpacket
		.response_empty         (adc_response_empty),              //               .empty
		.response_channel       (adc_response_channel),            //               .channel
		.response_data          (adc_response_data)                //               .data
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_adc_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
