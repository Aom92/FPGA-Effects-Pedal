-- REVERB.vhd

-- Generated using ACDS version 20.1 720

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity REVERB is
	port (
		ast_sink_data    : in  std_logic_vector(15 downto 0) := (others => '0'); --   avalon_streaming_sink.data
		ast_sink_valid   : in  std_logic                     := '0';             --                        .valid
		ast_sink_error   : in  std_logic_vector(1 downto 0)  := (others => '0'); --                        .error
		ast_source_data  : out std_logic_vector(46 downto 0);                    -- avalon_streaming_source.data
		ast_source_valid : out std_logic;                                        --                        .valid
		ast_source_error : out std_logic_vector(1 downto 0);                     --                        .error
		clk              : in  std_logic                     := '0';             --                     clk.clk
		reset_n          : in  std_logic                     := '0'              --                     rst.reset_n
	);
end entity REVERB;

architecture rtl of REVERB is
	component REVERB_fir_compiler_ii_0 is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset_n          : in  std_logic                     := 'X';             -- reset_n
			ast_sink_data    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			ast_sink_valid   : in  std_logic                     := 'X';             -- valid
			ast_sink_error   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			ast_source_data  : out std_logic_vector(46 downto 0);                    -- data
			ast_source_valid : out std_logic;                                        -- valid
			ast_source_error : out std_logic_vector(1 downto 0)                      -- error
		);
	end component REVERB_fir_compiler_ii_0;

begin

	fir_compiler_ii_0 : component REVERB_fir_compiler_ii_0
		port map (
			clk              => clk,              --                     clk.clk
			reset_n          => reset_n,          --                     rst.reset_n
			ast_sink_data    => ast_sink_data,    --   avalon_streaming_sink.data
			ast_sink_valid   => ast_sink_valid,   --                        .valid
			ast_sink_error   => ast_sink_error,   --                        .error
			ast_source_data  => ast_source_data,  -- avalon_streaming_source.data
			ast_source_valid => ast_source_valid, --                        .valid
			ast_source_error => ast_source_error  --                        .error
		);

end architecture rtl; -- of REVERB
