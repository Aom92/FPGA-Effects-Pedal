-- Effect_Pedal.vhd

-- Generated using ACDS version 20.1 720

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Effect_Pedal is
	port (
		adc_0_adc_response_valid         : out std_logic;                            -- adc_0_adc_response.valid
		adc_0_adc_response_startofpacket : out std_logic;                            --                   .startofpacket
		adc_0_adc_response_endofpacket   : out std_logic;                            --                   .endofpacket
		adc_0_adc_response_empty         : out std_logic_vector(0 downto 0);         --                   .empty
		adc_0_adc_response_channel       : out std_logic_vector(4 downto 0);         --                   .channel
		adc_0_adc_response_data          : out std_logic_vector(11 downto 0);        --                   .data
		adc_0_sample_clk_clk             : out std_logic;                            --   adc_0_sample_clk.clk
		clk_clk                          : in  std_logic                     := '0'; --                clk.clk
		reset_reset_n                    : in  std_logic                     := '0'  --              reset.reset_n
	);
end entity Effect_Pedal;

architecture rtl of Effect_Pedal is
	component Effect_Pedal_ADC_0 is
		port (
			adc_response_valid         : out std_logic;                            -- valid
			adc_response_startofpacket : out std_logic;                            -- startofpacket
			adc_response_endofpacket   : out std_logic;                            -- endofpacket
			adc_response_empty         : out std_logic_vector(0 downto 0);         -- empty
			adc_response_channel       : out std_logic_vector(4 downto 0);         -- channel
			adc_response_data          : out std_logic_vector(11 downto 0);        -- data
			clk_adc_clk                : in  std_logic                     := 'X'; -- clk
			reset_reset_n              : in  std_logic                     := 'X'; -- reset_n
			sample_clk_clk             : out std_logic                             -- clk
		);
	end component Effect_Pedal_ADC_0;

	component Effect_Pedal_Memory_Controller is
		port (
			clk_clk       : in std_logic := 'X'; -- clk
			reset_reset_n : in std_logic := 'X'  -- reset_n
		);
	end component Effect_Pedal_Memory_Controller;

begin

	adc_0 : component Effect_Pedal_ADC_0
		port map (
			adc_response_valid         => adc_0_adc_response_valid,         -- adc_response.valid
			adc_response_startofpacket => adc_0_adc_response_startofpacket, --             .startofpacket
			adc_response_endofpacket   => adc_0_adc_response_endofpacket,   --             .endofpacket
			adc_response_empty         => adc_0_adc_response_empty,         --             .empty
			adc_response_channel       => adc_0_adc_response_channel,       --             .channel
			adc_response_data          => adc_0_adc_response_data,          --             .data
			clk_adc_clk                => clk_clk,                          --      clk_adc.clk
			reset_reset_n              => reset_reset_n,                    --        reset.reset_n
			sample_clk_clk             => adc_0_sample_clk_clk              --   sample_clk.clk
		);

	memory_controller : component Effect_Pedal_Memory_Controller
		port map (
			clk_clk       => clk_clk,       --   clk.clk
			reset_reset_n => reset_reset_n  -- reset.reset_n
		);

end architecture rtl; -- of Effect_Pedal
