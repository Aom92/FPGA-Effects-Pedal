
module PWM_PLL (
	clk_clk,
	reset_reset_n,
	pwm_clk_clk);	

	input		clk_clk;
	input		reset_reset_n;
	output		pwm_clk_clk;
endmodule
